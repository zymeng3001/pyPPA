VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MACRO sky130_sram_0kbytes_1rw_32x512_32
   CLASS BLOCK ;
   SIZE 309.66 BY 899.78 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  107.08 0.0 107.46 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  112.92 0.0 113.3 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  118.76 0.0 119.14 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  124.6 0.0 124.98 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  130.44 0.0 130.82 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  136.28 0.0 136.66 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  142.12 0.0 142.5 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  147.96 0.0 148.34 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.8 0.0 154.18 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  159.64 0.0 160.02 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  165.48 0.0 165.86 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  171.32 0.0 171.7 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  177.16 0.0 177.54 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  183.0 0.0 183.38 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  188.84 0.0 189.22 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  194.68 0.0 195.06 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  200.52 0.0 200.9 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  206.36 0.0 206.74 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  212.2 0.0 212.58 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  218.04 0.0 218.42 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  223.88 0.0 224.26 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  229.72 0.0 230.1 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  235.56 0.0 235.94 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  247.24 0.0 247.62 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  253.08 0.0 253.46 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  258.92 0.0 259.3 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  264.76 0.0 265.14 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  270.6 0.0 270.98 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  276.44 0.0 276.82 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  282.28 0.0 282.66 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  288.12 0.0 288.5 0.38 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  293.96 0.0 294.34 0.38 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 137.17 0.38 137.55 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 145.67 0.38 146.05 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 151.31 0.38 151.69 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 159.81 0.38 160.19 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 165.45 0.38 165.83 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 173.95 0.38 174.33 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 179.59 0.38 179.97 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 188.09 0.38 188.47 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 193.585 0.38 193.965 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 201.985 0.38 202.365 ;
      END
   END addr0[9]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 14.87 0.38 15.25 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 23.37 0.38 23.75 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.1 0.0 31.48 0.38 ;
      END
   END clk0
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  299.8 0.0 300.18 0.38 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.045 0.0 179.425 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  183.69 0.0 184.07 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  185.425 0.0 185.805 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.515 0.0 186.895 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  189.53 0.0 189.91 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.835 0.0 193.215 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  195.425 0.0 195.805 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.895 0.0 198.275 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.715 0.0 199.095 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  202.895 0.0 203.275 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.045 0.0 204.425 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  207.895 0.0 208.275 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.045 0.0 209.425 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.895 0.0 213.275 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  214.045 0.0 214.425 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.73 0.0 219.11 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.425 0.0 220.805 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.075 0.0 222.455 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.57 0.0 224.95 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  227.895 0.0 228.275 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.425 0.0 230.805 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  232.895 0.0 233.275 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  233.755 0.0 234.135 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  237.895 0.0 238.275 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  239.045 0.0 239.425 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.895 0.0 243.275 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.045 0.0 244.425 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  247.93 0.0 248.31 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  249.045 0.0 249.425 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  253.77 0.0 254.15 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.425 0.0 255.805 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.115 0.0 257.495 0.38 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  259.61 0.0 259.99 0.38 ;
      END
   END dout0[32]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 309.04 899.16 ;
   LAYER  met2 ;
      RECT  0.62 0.62 309.04 899.16 ;
   LAYER  met3 ;
      RECT  0.98 0.62 309.04 136.57 ;
      RECT  0.98 136.57 309.04 138.15 ;
      RECT  0.98 138.15 309.04 899.16 ;
      RECT  0.62 138.15 0.98 145.07 ;
      RECT  0.62 146.65 0.98 150.71 ;
      RECT  0.62 152.29 0.98 159.21 ;
      RECT  0.62 160.79 0.98 164.85 ;
      RECT  0.62 166.43 0.98 173.35 ;
      RECT  0.62 174.93 0.98 178.99 ;
      RECT  0.62 180.57 0.98 187.49 ;
      RECT  0.62 189.07 0.98 192.985 ;
      RECT  0.62 194.565 0.98 201.385 ;
      RECT  0.62 202.965 0.98 899.16 ;
      RECT  0.62 0.62 0.98 14.27 ;
      RECT  0.62 15.85 0.98 22.77 ;
      RECT  0.62 24.35 0.98 136.57 ;
   LAYER  met4 ;
      RECT  0.62 0.98 106.48 899.16 ;
      RECT  106.48 0.98 108.06 899.16 ;
      RECT  108.06 0.98 309.04 899.16 ;
      RECT  108.06 0.62 112.32 0.98 ;
      RECT  113.9 0.62 118.16 0.98 ;
      RECT  119.74 0.62 124.0 0.98 ;
      RECT  125.58 0.62 129.84 0.98 ;
      RECT  131.42 0.62 135.68 0.98 ;
      RECT  137.26 0.62 141.52 0.98 ;
      RECT  143.1 0.62 147.36 0.98 ;
      RECT  148.94 0.62 153.2 0.98 ;
      RECT  154.78 0.62 159.04 0.98 ;
      RECT  160.62 0.62 164.88 0.98 ;
      RECT  166.46 0.62 170.72 0.98 ;
      RECT  172.3 0.62 176.56 0.98 ;
      RECT  265.74 0.62 270.0 0.98 ;
      RECT  271.58 0.62 275.84 0.98 ;
      RECT  277.42 0.62 281.68 0.98 ;
      RECT  283.26 0.62 287.52 0.98 ;
      RECT  289.1 0.62 293.36 0.98 ;
      RECT  0.62 0.62 30.5 0.98 ;
      RECT  32.08 0.62 106.48 0.98 ;
      RECT  294.94 0.62 299.2 0.98 ;
      RECT  300.78 0.62 309.04 0.98 ;
      RECT  178.14 0.62 178.445 0.98 ;
      RECT  180.025 0.62 182.4 0.98 ;
      RECT  184.67 0.62 184.825 0.98 ;
      RECT  187.495 0.62 188.24 0.98 ;
      RECT  190.51 0.62 192.235 0.98 ;
      RECT  193.815 0.62 194.08 0.98 ;
      RECT  196.405 0.62 197.295 0.98 ;
      RECT  199.695 0.62 199.92 0.98 ;
      RECT  201.5 0.62 202.295 0.98 ;
      RECT  205.025 0.62 205.76 0.98 ;
      RECT  210.025 0.62 211.6 0.98 ;
      RECT  215.025 0.62 217.44 0.98 ;
      RECT  219.71 0.62 219.825 0.98 ;
      RECT  221.405 0.62 221.475 0.98 ;
      RECT  223.055 0.62 223.28 0.98 ;
      RECT  225.55 0.62 227.295 0.98 ;
      RECT  228.875 0.62 229.12 0.98 ;
      RECT  231.405 0.62 232.295 0.98 ;
      RECT  234.735 0.62 234.96 0.98 ;
      RECT  236.54 0.62 237.295 0.98 ;
      RECT  240.025 0.62 240.8 0.98 ;
      RECT  245.025 0.62 246.64 0.98 ;
      RECT  250.025 0.62 252.48 0.98 ;
      RECT  254.75 0.62 254.825 0.98 ;
      RECT  256.405 0.62 256.515 0.98 ;
      RECT  258.095 0.62 258.32 0.98 ;
      RECT  260.59 0.62 264.16 0.98 ;
   END
END    sky130_sram_0kbytes_1rw_32x512_32
END    LIBRARY
