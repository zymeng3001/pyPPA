module chip_top (gpio);
	inout wire [63:0] gpio;
	wire clk;
	wire asyn_rst;
	wire IIN;
	wire EXT_CLK_IN;
	wire CLK_DIV_SEL_0;
	wire CLK_DIV_SEL_1;
	wire CLK_GATE_EN;
	wire CLK_DIV100;
	wire spi_clk;
	wire spi_csn;
	wire spi_mosi;
	wire spi_miso;
	wire qspi_clk;
	wire [15:0] qspi_mosi;
	wire qspi_mosi_valid;
	wire [15:0] qspi_miso;
	wire qspi_miso_valid;
	wire current_token_finish_flag;
	wire current_token_finish_work;
	wire qgen_state_work;
	wire qgen_state_end;
	wire kgen_state_work;
	wire kgen_state_end;
	wire vgen_state_work;
	wire vgen_state_end;
	wire att_qk_state_work;
	wire att_qk_state_end;
	wire att_pv_state_work;
	wire att_pv_state_end;
	wire proj_state_work;
	wire proj_state_end;
	wire ffn0_state_work;
	wire ffn0_state_end;
	wire ffn1_state_work;
	wire ffn1_state_end;
	CLK_GEN i_clk_gen(
		.asyn_rst(asyn_rst),
		.ext_clk(EXT_CLK_IN),
		.IIN(IIN),
		.clk_div_sel({CLK_DIV_SEL_1, CLK_DIV_SEL_0}),
		.clk_gate_en(CLK_GATE_EN),
		.o_chip_clk(clk),
		.o_clk_div(CLK_DIV100)
	);
	top top(
		.chip_clk(clk),
		.asyn_rst(asyn_rst),
		.spi_clk(spi_clk),
		.spi_csn(spi_csn),
		.spi_mosi(spi_mosi),
		.spi_miso(spi_miso),
		.qspi_clk(qspi_clk),
		.qspi_mosi(qspi_mosi),
		.qspi_mosi_valid(qspi_mosi_valid),
		.qspi_miso(qspi_miso),
		.qspi_miso_valid(qspi_miso_valid),
		.current_token_finish_flag(current_token_finish_flag),
		.current_token_finish_work(current_token_finish_work),
		.qgen_state_work(qgen_state_work),
		.qgen_state_end(qgen_state_end),
		.kgen_state_work(kgen_state_work),
		.kgen_state_end(kgen_state_end),
		.vgen_state_work(vgen_state_work),
		.vgen_state_end(vgen_state_end),
		.att_qk_state_work(att_qk_state_work),
		.att_qk_state_end(att_qk_state_end),
		.att_pv_state_work(att_pv_state_work),
		.att_pv_state_end(att_pv_state_end),
		.proj_state_work(proj_state_work),
		.proj_state_end(proj_state_end),
		.ffn0_state_work(ffn0_state_work),
		.ffn0_state_end(ffn0_state_end),
		.ffn1_state_work(ffn1_state_work),
		.ffn1_state_end(ffn1_state_end)
	);
	sdio_1v8_n1 south_io_0(
		.outi(asyn_rst),
		.outi_1v8(),
		.pad(gpio[0]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_1(
		.outi(spi_clk),
		.outi_1v8(),
		.pad(gpio[1]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_2(
		.outi(spi_csn),
		.outi_1v8(),
		.pad(gpio[2]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_3(
		.outi(spi_mosi),
		.outi_1v8(),
		.pad(gpio[3]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_4(
		.outi(),
		.outi_1v8(),
		.pad(gpio[4]),
		.ana_io_1v8(),
		.dq(~spi_miso),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_5(
		.outi(qspi_clk),
		.outi_1v8(),
		.pad(gpio[5]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_6(
		.outi(qspi_mosi[0]),
		.outi_1v8(),
		.pad(gpio[6]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_7(
		.outi(qspi_mosi[1]),
		.outi_1v8(),
		.pad(gpio[7]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_8(
		.outi(qspi_mosi[2]),
		.outi_1v8(),
		.pad(gpio[8]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_9(
		.outi(qspi_mosi[3]),
		.outi_1v8(),
		.pad(gpio[9]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_10(
		.outi(qspi_mosi[4]),
		.outi_1v8(),
		.pad(gpio[10]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_11(
		.outi(qspi_mosi[5]),
		.outi_1v8(),
		.pad(gpio[11]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_12(
		.outi(qspi_mosi[6]),
		.outi_1v8(),
		.pad(gpio[12]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_13(
		.outi(qspi_mosi[7]),
		.outi_1v8(),
		.pad(gpio[13]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_14(
		.outi(qspi_mosi[8]),
		.outi_1v8(),
		.pad(gpio[14]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_15(
		.outi(qspi_mosi[9]),
		.outi_1v8(),
		.pad(gpio[15]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_16(
		.outi(qspi_mosi[10]),
		.outi_1v8(),
		.pad(gpio[16]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_17(
		.outi(qspi_mosi[11]),
		.outi_1v8(),
		.pad(gpio[17]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_18(
		.outi(qspi_mosi[12]),
		.outi_1v8(),
		.pad(gpio[18]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_19(
		.outi(qspi_mosi[13]),
		.outi_1v8(),
		.pad(gpio[19]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_20(
		.outi(qspi_mosi[14]),
		.outi_1v8(),
		.pad(gpio[20]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_21(
		.outi(qspi_mosi[15]),
		.outi_1v8(),
		.pad(gpio[21]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_22(
		.outi(qspi_mosi_valid),
		.outi_1v8(),
		.pad(gpio[22]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_23(
		.outi(),
		.outi_1v8(),
		.pad(gpio[23]),
		.ana_io_1v8(),
		.dq(~qspi_miso[0]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_24(
		.outi(),
		.outi_1v8(),
		.pad(gpio[24]),
		.ana_io_1v8(),
		.dq(~qspi_miso[1]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_25(
		.outi(),
		.outi_1v8(),
		.pad(gpio[25]),
		.ana_io_1v8(),
		.dq(~qspi_miso[2]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_26(
		.outi(),
		.outi_1v8(),
		.pad(gpio[26]),
		.ana_io_1v8(),
		.dq(~qspi_miso[3]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_27(
		.outi(),
		.outi_1v8(),
		.pad(gpio[27]),
		.ana_io_1v8(),
		.dq(~qspi_miso[4]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_28(
		.outi(),
		.outi_1v8(),
		.pad(gpio[28]),
		.ana_io_1v8(),
		.dq(~qspi_miso[5]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_29(
		.outi(),
		.outi_1v8(),
		.pad(gpio[29]),
		.ana_io_1v8(),
		.dq(~qspi_miso[6]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_30(
		.outi(),
		.outi_1v8(),
		.pad(gpio[30]),
		.ana_io_1v8(),
		.dq(~qspi_miso[7]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_31(
		.outi(),
		.outi_1v8(),
		.pad(gpio[31]),
		.ana_io_1v8(),
		.dq(~qspi_miso[8]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_32(
		.outi(),
		.outi_1v8(),
		.pad(gpio[32]),
		.ana_io_1v8(),
		.dq(~qspi_miso[9]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_33(
		.outi(),
		.outi_1v8(),
		.pad(gpio[33]),
		.ana_io_1v8(),
		.dq(~qspi_miso[10]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_34(
		.outi(),
		.outi_1v8(),
		.pad(gpio[34]),
		.ana_io_1v8(),
		.dq(~qspi_miso[11]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_35(
		.outi(),
		.outi_1v8(),
		.pad(gpio[35]),
		.ana_io_1v8(),
		.dq(~qspi_miso[12]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_36(
		.outi(),
		.outi_1v8(),
		.pad(gpio[36]),
		.ana_io_1v8(),
		.dq(~qspi_miso[13]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_37(
		.outi(),
		.outi_1v8(),
		.pad(gpio[37]),
		.ana_io_1v8(),
		.dq(~qspi_miso[14]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_38(
		.outi(),
		.outi_1v8(),
		.pad(gpio[38]),
		.ana_io_1v8(),
		.dq(~qspi_miso[15]),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 south_io_39(
		.outi(),
		.outi_1v8(),
		.pad(gpio[39]),
		.ana_io_1v8(),
		.dq(~qspi_miso_valid),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_1(
		.outi(EXT_CLK_IN),
		.outi_1v8(),
		.pad(gpio[41]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_2(
		.outi(CLK_DIV_SEL_0),
		.outi_1v8(),
		.pad(gpio[42]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_3(
		.outi(CLK_DIV_SEL_1),
		.outi_1v8(),
		.pad(gpio[43]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_4(
		.outi(CLK_GATE_EN),
		.outi_1v8(),
		.pad(gpio[44]),
		.ana_io_1v8(),
		.dq(1'b0),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b1),
		.pd(1'b1),
		.ppen(1'b0),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_5(
		.outi(),
		.outi_1v8(),
		.pad(gpio[45]),
		.ana_io_1v8(),
		.dq(~CLK_DIV100),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_6(
		.outi(),
		.outi_1v8(),
		.pad(gpio[46]),
		.ana_io_1v8(),
		.dq(~current_token_finish_flag),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_7(
		.outi(),
		.outi_1v8(),
		.pad(gpio[47]),
		.ana_io_1v8(),
		.dq(~current_token_finish_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_8(
		.outi(),
		.outi_1v8(),
		.pad(gpio[48]),
		.ana_io_1v8(),
		.dq(~qgen_state_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_9(
		.outi(),
		.outi_1v8(),
		.pad(gpio[49]),
		.ana_io_1v8(),
		.dq(~qgen_state_end),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_10(
		.outi(),
		.outi_1v8(),
		.pad(gpio[50]),
		.ana_io_1v8(),
		.dq(~kgen_state_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_11(
		.outi(),
		.outi_1v8(),
		.pad(gpio[51]),
		.ana_io_1v8(),
		.dq(~kgen_state_end),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_12(
		.outi(),
		.outi_1v8(),
		.pad(gpio[52]),
		.ana_io_1v8(),
		.dq(~vgen_state_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_13(
		.outi(),
		.outi_1v8(),
		.pad(gpio[53]),
		.ana_io_1v8(),
		.dq(~vgen_state_end),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_14(
		.outi(),
		.outi_1v8(),
		.pad(gpio[54]),
		.ana_io_1v8(),
		.dq(~att_qk_state_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_15(
		.outi(),
		.outi_1v8(),
		.pad(gpio[55]),
		.ana_io_1v8(),
		.dq(~att_qk_state_end),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_16(
		.outi(),
		.outi_1v8(),
		.pad(gpio[56]),
		.ana_io_1v8(),
		.dq(~att_pv_state_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_17(
		.outi(),
		.outi_1v8(),
		.pad(gpio[57]),
		.ana_io_1v8(),
		.dq(~att_pv_state_end),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_18(
		.outi(),
		.outi_1v8(),
		.pad(gpio[58]),
		.ana_io_1v8(),
		.dq(~proj_state_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_19(
		.outi(),
		.outi_1v8(),
		.pad(gpio[59]),
		.ana_io_1v8(),
		.dq(~proj_state_end),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_20(
		.outi(),
		.outi_1v8(),
		.pad(gpio[60]),
		.ana_io_1v8(),
		.dq(~ffn0_state_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_21(
		.outi(),
		.outi_1v8(),
		.pad(gpio[61]),
		.ana_io_1v8(),
		.dq(~ffn0_state_end),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_22(
		.outi(),
		.outi_1v8(),
		.pad(gpio[62]),
		.ana_io_1v8(),
		.dq(~ffn1_state_work),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
	sdio_1v8_n1 north_io_23(
		.outi(),
		.outi_1v8(),
		.pad(gpio[63]),
		.ana_io_1v8(),
		.dq(~ffn1_state_end),
		.drv0(1'b0),
		.drv1(1'b0),
		.drv2(1'b0),
		.enabq(1'b0),
		.enq(1'b0),
		.pd(1'b1),
		.ppen(1'b1),
		.prg_slew(1'b0),
		.puq(1'b1),
		.pwrupzhl(1'b0),
		.pwrup_pull_en(1'b0)
	);
endmodule
